library ieee;
use ieee.std_logic_1164.all;

entity datapath is
	port(
		constant_in : in STD_LOGIC_VECTOR (15 downto 0);
        MB_select : in STD_LOGIC;
        MD_select : in STD_LOGIC;
        data_in : in STD_LOGIC_VECTOR (15 downto 0);
        clk : in STD_LOGIC;
        write : in STD_LOGIC;
        D_address : in STD_LOGIC_VECTOR(2 downto 0);
        A_address : in STD_LOGIC_VECTOR(2 downto 0);
        B_address : in STD_LOGIC_VECTOR(2 downto 0);
        FS : in STD_LOGIC_VECTOR(4 downto 0);
        address_out : out STD_LOGIC_VECTOR (15 downto 0);
        data_out : out STD_LOGIC_VECTOR (15 downto 0);
        V : out STD_LOGIC;
        C : out STD_LOGIC;
        N : out STD_LOGIC;
        Z : out STD_LOGIC);
end datapath;

architecture behavioral of datapath is

	component register_file port(
		load_enable : in STD_LOGIC;
		clk : in STD_LOGIC;
		data : in STD_LOGIC_VECTOR(15 downto 0);
		A_select : in STD_LOGIC_VECTOR(2 downto 0);
		B_select : in STD_LOGIC_VECTOR(2 downto 0);
		D_select : in STD_LOGIC_VECTOR(2 downto 0);
		A_data : out STD_LOGIC_VECTOR(15 downto 0);
		B_data : out STD_LOGIC_VECTOR(15 downto 0));
	end component;

	component function_unit port(
		A : in std_logic_vector (15 downto 0);
        B : in std_logic_vector (15 downto 0);
        FS : in std_logic_vector (4 downto 0);
		V : out std_logic;
		C : out std_logic;
		N : out std_logic;
		Z : out std_logic;
		F : out std_logic_vector (15 downto 0));
	end component;

	component mux2_16 port(
		in0 : in STD_LOGIC_VECTOR (15 downto 0);
		in1 : in STD_LOGIC_VECTOR (15 downto 0);
		S : in STD_LOGIC;
		Z : out STD_LOGIC_VECTOR (15 downto 0));
	end component;

	signal functional_unit_out : STD_LOGIC_VECTOR(15 downto 0);
	signal muxB_out : STD_LOGIC_VECTOR(15 downto 0);
	signal muxD_out : STD_LOGIC_VECTOR(15 downto 0);
	signal A_data_out : STD_LOGIC_VECTOR(15 downto 0);
	signal B_data_out : STD_LOGIC_VECTOR(15 downto 0);

begin

	function_unit : function_unit port map(
		A=>A_data_out,
		B=>muxB_out,
		FS=>FS,
		F=>functional_unit_out,
		V=>V,
		C=>C,
		N=>N,
		Z=>Z);

	muxB : mux2_16 port map(
		in0 => B_data_out,
		in1 => constant_in,
		S => MB_select,
		Z => muxB_out);

	muxD : mux2_16 port map(
		in0 => functional_unit_out,
		in1 => data_in,
		S => MD_select,
		Z => muxD_out);

end behavioral;
