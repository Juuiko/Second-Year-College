library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity reg4 is
	port(
		D : in std_logic_vector(3 downto 0);
		load : in std_logic;
		Clk : in std_logic;
		Q : out std_logic_vector(3 downto 0));
end reg4;

architecture Behavioral of reg4 is
begin
	process(Clk)
	begin
		if (rising_edge(Clk)) then
			if load='1' then
				Q<=D after 5 ns;
			end if;
		end if;
	end process;
end Behavioral;
